`timescale 1ns / 1ps


module VGA_Controller (
    input  logic clk,         // 시스템 클럭 (예: 100MHz)
    input  logic reset,       // 비동기 리셋
    output logic rclk,
    output logic h_sync,      // VGA HSync
    output logic v_sync,      // VGA VSync
    output logic [9:0] x_pixel, // 현재 유효 픽셀의 x 좌표
    output logic [9:0] y_pixel, // 현재 유효 픽셀의 y 좌표
    output logic DE,
    output logic pclk          // Display Enable (유효 픽셀 출력 여부)
);

    // 내부 신호
    logic [9:0]  h_counter;
    logic [9:0]  v_counter;

    assign rclk = clk;

    // 1. 픽셀 클럭 생성기 인스턴스
    pixel_clk_gen u_clk_gen (
        .clk     (clk),
        .reset   (reset),
        .pclk    (pclk)
    );

    // 2. 픽셀 카운터 인스턴스
    pixel_counter u_counter (
        .pclk      (pclk),
        .reset     (reset),
        .h_counter (h_counter),
        .v_counter (v_counter)
    );

    // 3. VGA 타이밍 디코더 인스턴스
    vga_decoder u_decoder (
        .h_counter (h_counter),
        .v_counter (v_counter),
        .h_sync    (h_sync),
        .v_sync    (v_sync),
        .x_pixel   (x_pixel),
        .y_pixel   (y_pixel),
        .DE        (DE)
    );

endmodule






module pixel_clk_gen (
    input logic clk,
    input logic reset,
    output logic pclk
);

    logic [1:0] p_counter;

    always_ff @( posedge clk or posedge reset ) begin 
        if (reset) begin
            p_counter <=0;
            pclk <=0;
        end else begin
            if (p_counter == 4-1) begin
                p_counter <= 0;
                pclk <= 1;
            end else begin
                p_counter <= p_counter+1;
                pclk <= 0;
            end
        end
    end


    
endmodule


module pixel_counter (
    input logic pclk,
    input logic reset,
    output logic [9:0] h_counter,
    output logic [9:0] v_counter
);

    localparam H_MAX = 800, V_MAX = 525;

    // Horizontal Count    
    always_ff @( posedge pclk or posedge reset ) begin 
        if (reset) begin
            h_counter <=0;
        end else begin
            if (h_counter == H_MAX -1) begin
                h_counter <= 0;
            end else begin
                h_counter <= h_counter + 1;
            end
        end
        
    end

    // Vertical Count
    always_ff @( posedge pclk or posedge reset ) begin : blockName
        if (reset) begin
            v_counter <= 0;
        end else begin
            if (h_counter == H_MAX -1) begin
                if (v_counter == V_MAX -1 ) begin
                    v_counter <= 0;
                end else begin
                    v_counter <= v_counter+1;
                end
            end
        end
    end


endmodule



module vga_decoder (
    input logic [9:0] h_counter,
    input logic [9:0] v_counter,
    output logic h_sync,
    output logic v_sync,
    output logic [9:0] x_pixel,
    output logic [9:0] y_pixel,
    output logic DE
);
    

    localparam H_Visible_area	=640;
    localparam H_Front_porch	=16;	
    localparam H_Sync_pulse	=96;
    localparam H_Back_porch	=48;	
    localparam H_Whole_line	=800;	

    localparam V_Visible_area	=480;	
    localparam V_Front_porch	=10;	
    localparam V_Sync_pulse	=2;	
    localparam V_Back_porch	=33;	
    localparam V_Whole_frame =525;	


    assign h_sync = !((h_counter >= (H_Visible_area + H_Front_porch)) &&
                    (h_counter < (H_Visible_area + H_Front_porch + H_Sync_pulse)) );


    assign v_sync = !((v_counter >= (V_Visible_area + V_Front_porch)) &&
                    (v_counter < (V_Visible_area + V_Front_porch + V_Sync_pulse)) );


    assign DE = (h_counter < H_Visible_area) && (v_counter < V_Visible_area);


    assign x_pixel = h_counter;
    assign y_pixel = v_counter;  

endmodule