`timescale 1ns / 1ps
module rom_command(
    input  logic [7:0] char_code,
    input  logic [3:0] row,        // 0~15
    output logic [15:0] font_bits
);

    logic [15:0] rom [0:127][0:15];

    initial begin
        // W
        rom["W"][0]  = 16'b1100000000000011;
        rom["W"][1]  = 16'b1100000000000011;
        rom["W"][2]  = 16'b1100000000000011;
        rom["W"][3]  = 16'b1100000000000011;
        rom["W"][4]  = 16'b1100000000000011;
        rom["W"][5]  = 16'b1100000000000011;
        rom["W"][6]  = 16'b1100001100000011;
        rom["W"][7]  = 16'b1100001100000011;
        rom["W"][8]  = 16'b1100001100000011;
        rom["W"][9]  = 16'b1100001100000011;
        rom["W"][10] = 16'b0110011001100110;
        rom["W"][11] = 16'b0110011001100110;
        rom["W"][12] = 16'b0011110001111100;
        rom["W"][13] = 16'b0011110001111100;
        rom["W"][14] = 16'b0000000000000000;
        rom["W"][15] = 16'b0000000000000000;

        // A
        rom["A"][0]  = 16'b0000001100000000;
        rom["A"][1]  = 16'b0000011110000000;
        rom["A"][2]  = 16'b0000110011000000;
        rom["A"][3]  = 16'b0001100001100000;
        rom["A"][4]  = 16'b0001100001100000;
        rom["A"][5]  = 16'b0011000000110000;
        rom["A"][6]  = 16'b0011111111110000;
        rom["A"][7]  = 16'b0011111111110000;
        rom["A"][8]  = 16'b0110000000011000;
        rom["A"][9]  = 16'b0110000000011000;
        rom["A"][10] = 16'b1100000000001100;
        rom["A"][11] = 16'b1100000000001100;
        rom["A"][12] = 16'b1100000000001100;
        rom["A"][13] = 16'b0000000000000000;
        rom["A"][14] = 16'b0000000000000000;
        rom["A"][15] = 16'b0000000000000000;

        // R
        rom["R"][0]  = 16'b0111111111100000;
        rom["R"][1]  = 16'b0111111111110000;
        rom["R"][2]  = 16'b0011000000110000;
        rom["R"][3]  = 16'b0011000000110000;
        rom["R"][4]  = 16'b0011000000110000;
        rom["R"][5]  = 16'b0011111111110000;
        rom["R"][6]  = 16'b0011111111100000;
        rom["R"][7]  = 16'b0011000111000000;
        rom["R"][8]  = 16'b0011000011000000;
        rom["R"][9]  = 16'b0011000011100000;
        rom["R"][10] = 16'b0011000001110000;
        rom["R"][11] = 16'b0011000000110000;
        rom["R"][12] = 16'b0000000000000000;
        rom["R"][13] = 16'b0000000000000000;
        rom["R"][14] = 16'b0000000000000000;
        rom["R"][15] = 16'b0000000000000000;

        // N
        rom["N"][0]  = 16'b1100000000110000;
        rom["N"][1]  = 16'b1110000000110000;
        rom["N"][2]  = 16'b1011000000110000;
        rom["N"][3]  = 16'b1001100000110000;
        rom["N"][4]  = 16'b1000110000110000;
        rom["N"][5]  = 16'b1000011000110000;
        rom["N"][6]  = 16'b1000001100110000;
        rom["N"][7]  = 16'b1000000110110000;
        rom["N"][8]  = 16'b1000000011110000;
        rom["N"][9]  = 16'b1000000001110000;
        rom["N"][10] = 16'b1000000000110000;
        rom["N"][11] = 16'b1000000000110000;
        rom["N"][12] = 16'b0000000000000000;
        rom["N"][13] = 16'b0000000000000000;
        rom["N"][14] = 16'b0000000000000000;
        rom["N"][15] = 16'b0000000000000000;

        // I
        rom["I"][0]  = 16'b0001111111100000;
        rom["I"][1]  = 16'b0000011000000000;
        rom["I"][2]  = 16'b0000011000000000;
        rom["I"][3]  = 16'b0000011000000000;
        rom["I"][4]  = 16'b0000011000000000;
        rom["I"][5]  = 16'b0000011000000000;
        rom["I"][6]  = 16'b0000011000000000;
        rom["I"][7]  = 16'b0000011000000000;
        rom["I"][8]  = 16'b0000011000000000;
        rom["I"][9]  = 16'b0000011000000000;
        rom["I"][10] = 16'b0001111111100000;
        rom["I"][11] = 16'b0000000000000000;
        rom["I"][12] = 16'b0000000000000000;
        rom["I"][13] = 16'b0000000000000000;
        rom["I"][14] = 16'b0000000000000000;
        rom["I"][15] = 16'b0000000000000000;

        // G
        rom["G"][0]  = 16'b0001111111100000;
        rom["G"][1]  = 16'b0011000000110000;
        rom["G"][2]  = 16'b0110000000000000;
        rom["G"][3]  = 16'b0110000000000000;
        rom["G"][4]  = 16'b0110001111110000;
        rom["G"][5]  = 16'b0110000000110000;
        rom["G"][6]  = 16'b0110000000110000;
        rom["G"][7]  = 16'b0110000000110000;
        rom["G"][8]  = 16'b0011000000110000;
        rom["G"][9]  = 16'b0001111111100000;
        rom["G"][10] = 16'b0000000000000000;
        rom["G"][11] = 16'b0000000000000000;
        rom["G"][12] = 16'b0000000000000000;
        rom["G"][13] = 16'b0000000000000000;
        rom["G"][14] = 16'b0000000000000000;
        rom["G"][15] = 16'b0000000000000000;
    end

    assign font_bits = rom[char_code][row];
endmodule
